LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY codificador IS PORT (
	s: IN STD_LOGIC_VECTOR(0 to 7);
	o: OUT STD_LOGIC_VECTOR(2 downto 0)
	);
END codificador;

ARCHITECTURE arq OF codificador IS

BEGIN
	WITH s SELECT
		o <= 
			"000" WHEN "10000000",
			"001" WHEN "01000000",
			"010" WHEN "00100000",
			"011" WHEN "00010000",
			"100" WHEN "00001000",
			"101" WHEN "00000100",
			"110" WHEN "00000010",
			"111" WHEN "00000001",
			"000" WHEN OTHERS;		
END arq;