LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY demux1x4 IS PORT (
	f: IN STD_LOGIC;
	x : OUT STD_LOGIC_VECTOR(3 downto 0);
	s: IN STD_LOGIC_VECTOR(1 downto 0)
	);
END demux1x4;

ARCHITECTURE demux OF demux1x4 IS

BEGIN
	WITH s SELECT
		x(0) <= f WHEN "00", '0' WHEN OTHERS;
		
	WITH s SELECT
		x(1) <= f WHEN "01", '0' WHEN OTHERS;

	WITH s SELECT
		x(2) <= f WHEN "10", '0' WHEN OTHERS;
		
	WITH s SELECT
		x(3) <= f WHEN "11", '0' WHEN OTHERS;
END demux;
	